reg [19:0] C_LATCH;
reg [15:0] S_LATCH;

assign {46,45,44,43,41,40,39,38,14,13,12,11,9,8,7,6,33,32,1,64} = C_LATCH;
assign {37,36,35,34,18,17,16,15,5,4,3,2,51,50,49,48} = S_LATCH;
assign 47 = ~46;

always @(posedge 23)
  C_LATCH <= {27,25,59,57,55,54,53,52,31,30,29,28,22,21,20,19,63,62,61,60};

always @(posedge 24)
  S_LATCH <= {55,54,53,52,31,30,29,28,22,21,20,19,63,62,61,60};
